`timescale 1ns/1ps

module hsv2rgb(
    input      [6:0]     i_hsv,
    output reg [23:0]    o_rgb
);

always @ (*) begin
    case (i_hsv)
    //                  rrggbb //NESDoc.pdf
    7'h00:  o_rgb = 24'h757575;//24'h000000;
    7'h01:  o_rgb = 24'h271B8F;//24'h000000;
    7'h02:  o_rgb = 24'h0000AB;//24'h000000;
    7'h03:  o_rgb = 24'h47009F;//24'h000000;
    7'h04:  o_rgb = 24'h8F0077;//24'h000000;
    7'h05:  o_rgb = 24'hAB0013;//24'h000000;
    7'h06:  o_rgb = 24'hA70000;//24'h000000;
    7'h07:  o_rgb = 24'h7F0B00;//24'h000000;
    7'h08:  o_rgb = 24'h432F00;//24'h000000;
    7'h09:  o_rgb = 24'h004700;//24'h000000;
    7'h0A:  o_rgb = 24'h005100;//24'h000000;
    7'h0B:  o_rgb = 24'h003F17;//24'h000000;
    7'h0C:  o_rgb = 24'h1B3F5F;//24'h000000;
    7'h0D:  o_rgb = 24'h000000;//24'h000000;
    7'h0E:  o_rgb = 24'h000000;//24'h000000;
    7'h0F:  o_rgb = 24'h000000;//24'h000000;
    7'h10:  o_rgb = 24'hBCBCBC;//24'h404040;
    7'h11:  o_rgb = 24'h0073EF;//24'h404040;
    7'h12:  o_rgb = 24'h233BEF;//24'h404040;
    7'h13:  o_rgb = 24'h8300F3;//24'h404040;
    7'h14:  o_rgb = 24'hBF00BF;//24'h404040;
    7'h15:  o_rgb = 24'hE7005B;//24'h404040;
    7'h16:  o_rgb = 24'hDB2B00;//24'h404040;
    7'h17:  o_rgb = 24'hCB4F0F;//24'h404040;
    7'h18:  o_rgb = 24'h8B7300;//24'h404040;
    7'h19:  o_rgb = 24'h009700;//24'h404040;
    7'h1A:  o_rgb = 24'h00AB00;//24'h404040;
    7'h1B:  o_rgb = 24'h00933B;//24'h404040;
    7'h1C:  o_rgb = 24'h00838B;//24'h404040;
    7'h1D:  o_rgb = 24'h000000;//24'h404040;
    7'h1E:  o_rgb = 24'h000000;//24'h404040;
    7'h1F:  o_rgb = 24'h000000;//24'h404040;
    7'h20:  o_rgb = 24'hFFFFFF;//24'h808080;
    7'h21:  o_rgb = 24'h3FBFFF;//24'h808080;
    7'h22:  o_rgb = 24'h5F97FF;//24'h808080;
    7'h23:  o_rgb = 24'hA78BFD;//24'h808080;
    7'h24:  o_rgb = 24'hF77BFF;//24'h808080;
    7'h25:  o_rgb = 24'hFF77B7;//24'h808080;
    7'h26:  o_rgb = 24'hFF7763;//24'h808080;
    7'h27:  o_rgb = 24'hFF9B3B;//24'h808080;
    7'h28:  o_rgb = 24'hF3BF3F;//24'h808080;
    7'h29:  o_rgb = 24'h83D313;//24'h808080;
    7'h2A:  o_rgb = 24'h4FDF4B;//24'h808080;
    7'h2B:  o_rgb = 24'h58F898;//24'h808080;
    7'h2C:  o_rgb = 24'h00EBDB;//24'h808080;
    7'h2D:  o_rgb = 24'h000000;//24'h808080;
    7'h2E:  o_rgb = 24'h000000;//24'h808080;
    7'h2F:  o_rgb = 24'h000000;//24'h808080;
    7'h30:  o_rgb = 24'hFFFFFF;//24'hc0c0c0;
    7'h31:  o_rgb = 24'hABE7FF;//24'hc0c0c0;
    7'h32:  o_rgb = 24'hC7D7FF;//24'hc0c0c0;
    7'h33:  o_rgb = 24'hD7CBFF;//24'hc0c0c0;
    7'h34:  o_rgb = 24'hFFC7FF;//24'hc0c0c0;
    7'h35:  o_rgb = 24'hFFC7DB;//24'hc0c0c0;
    7'h36:  o_rgb = 24'hFFBFB3;//24'hc0c0c0;
    7'h37:  o_rgb = 24'hFFDBAB;//24'hc0c0c0;
    7'h38:  o_rgb = 24'hFFE7A3;//24'hc0c0c0;
    7'h39:  o_rgb = 24'hE3FFA3;//24'hc0c0c0;
    7'h3A:  o_rgb = 24'hABF3BF;//24'hc0c0c0;
    7'h3B:  o_rgb = 24'hB3FFCF;//24'hc0c0c0;
    7'h3C:  o_rgb = 24'h9FFFF3;//24'hc0c0c0;
    7'h3D:  o_rgb = 24'h000000;//24'hc0c0c0;
    7'h3E:  o_rgb = 24'h000000;//24'hc0c0c0;
    7'h3F:  o_rgb = 24'h000000;//24'hc0c0c0;
    7'h40:  o_rgb = 24'h757575;//24'h000000;
    7'h41:  o_rgb = 24'h271B8F;//24'h000000;
    7'h42:  o_rgb = 24'h0000AB;//24'h000000;
    7'h43:  o_rgb = 24'h47009F;//24'h000000;
    7'h44:  o_rgb = 24'h8F0077;//24'h000000;
    7'h45:  o_rgb = 24'hAB0013;//24'h000000;
    7'h46:  o_rgb = 24'hA70000;//24'h000000;
    7'h47:  o_rgb = 24'h7F0B00;//24'h000000;
    7'h48:  o_rgb = 24'h432F00;//24'h000000;
    7'h49:  o_rgb = 24'h004700;//24'h000000;
    7'h4A:  o_rgb = 24'h005100;//24'h000000;
    7'h4B:  o_rgb = 24'h003F17;//24'h000000;
    7'h4C:  o_rgb = 24'h1B3F5F;//24'h000000;
    7'h4D:  o_rgb = 24'h000000;//24'h000000;
    7'h4E:  o_rgb = 24'h000000;//24'h000000;
    7'h4F:  o_rgb = 24'h000000;//24'h000000;
    7'h50:  o_rgb = 24'hBCBCBC;//24'h400000;
    7'h51:  o_rgb = 24'h0073EF;//24'h401800;
    7'h52:  o_rgb = 24'h233BEF;//24'h403000;
    7'h53:  o_rgb = 24'h8300F3;//24'h384000;
    7'h54:  o_rgb = 24'hBF00BF;//24'h204000;
    7'h55:  o_rgb = 24'hE7005B;//24'h084000;
    7'h56:  o_rgb = 24'hDB2B00;//24'h004010;
    7'h57:  o_rgb = 24'hCB4F0F;//24'h004028;
    7'h58:  o_rgb = 24'h8B7300;//24'h004040;
    7'h59:  o_rgb = 24'h009700;//24'h002840;
    7'h5A:  o_rgb = 24'h00AB00;//24'h001040;
    7'h5B:  o_rgb = 24'h00933B;//24'h080040;
    7'h5C:  o_rgb = 24'h00838B;//24'h200040;
    7'h5D:  o_rgb = 24'h000000;//24'h380040;
    7'h5E:  o_rgb = 24'h000000;//24'h400030;
    7'h5F:  o_rgb = 24'h000000;//24'h400018;
    7'h60:  o_rgb = 24'hFFFFFF;//24'h800000;
    7'h61:  o_rgb = 24'h3FBFFF;//24'h803000;
    7'h62:  o_rgb = 24'h5F97FF;//24'h806000;
    7'h63:  o_rgb = 24'hA78BFD;//24'h708000;
    7'h64:  o_rgb = 24'hF77BFF;//24'h408000;
    7'h65:  o_rgb = 24'hFF77B7;//24'h108000;
    7'h66:  o_rgb = 24'hFF7763;//24'h008020;
    7'h67:  o_rgb = 24'hFF9B3B;//24'h008050;
    7'h68:  o_rgb = 24'hF3BF3F;//24'h008080;
    7'h69:  o_rgb = 24'h83D313;//24'h005080;
    7'h6A:  o_rgb = 24'h4FDF4B;//24'h002080;
    7'h6B:  o_rgb = 24'h58F898;//24'h100080;
    7'h6C:  o_rgb = 24'h00EBDB;//24'h400080;
    7'h6D:  o_rgb = 24'h000000;//24'h700080;
    7'h6E:  o_rgb = 24'h000000;//24'h800060;
    7'h6F:  o_rgb = 24'h000000;//24'h800030;
    7'h70:  o_rgb = 24'hFFFFFF;//24'hc00000;
    7'h71:  o_rgb = 24'hABE7FF;//24'hc04800;
    7'h72:  o_rgb = 24'hC7D7FF;//24'hc09000;
    7'h73:  o_rgb = 24'hD7CBFF;//24'ha8c000;
    7'h74:  o_rgb = 24'hFFC7FF;//24'h60c000;
    7'h75:  o_rgb = 24'hFFC7DB;//24'h18c000;
    7'h76:  o_rgb = 24'hFFBFB3;//24'h00c030;
    7'h77:  o_rgb = 24'hFFDBAB;//24'h00c078;
    7'h78:  o_rgb = 24'hFFE7A3;//24'h00c0c0;
    7'h79:  o_rgb = 24'hE3FFA3;//24'h0078c0;
    7'h7A:  o_rgb = 24'hABF3BF;//24'h0030c0;
    7'h7B:  o_rgb = 24'hB3FFCF;//24'h1800c0;
    7'h7C:  o_rgb = 24'h9FFFF3;//24'h6000c0;
    7'h7D:  o_rgb = 24'h000000;//24'ha800c0;
    7'h7E:  o_rgb = 24'h000000;//24'hc00090;
    7'h7F:  o_rgb = 24'h000000;//24'hc00048;
    endcase
end
endmodule
module ppu_rde(
);

endmodule
